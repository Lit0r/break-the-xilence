--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   07:23:48 01/07/2014
-- Design Name:   
-- Module Name:   C:/Users/hamster/Projects/FPGA/adau1761_test/tb_adau1761_test.vhd
-- Project Name:  adau1761_test
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: adau1761_test
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types- always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
ENTITY tb_adau1761_test IS
END tb_adau1761_test;
 
ARCHITECTURE behavior OF tb_adau1761_test IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
	COMPONENT adau1761_test
	PORT(
		clk_100 : IN std_logic;
		AC_GPIO1 : IN std_logic;
		AC_GPIO2 : IN std_logic;
		AC_GPIO3 : IN std_logic;    
		AC_SDA : INOUT std_logic;      
		AC_ADR0 : OUT std_logic;
		AC_ADR1 : OUT std_logic;
		AC_GPIO0 : OUT std_logic;
		AC_MCLK : OUT std_logic;
		AC_SCK : OUT std_logic;
           sw       : in    STD_LOGIC_VECTOR(7 downto 0)
           
		);
	END COMPONENT;    

   --Inputs
   signal clk_100 : std_logic := '0';
   signal AC_GPIO1 : std_logic := '0';

	--BiDirs
   signal AC_SDA : std_logic;

 	--Outputs
   signal AC_ADR0 : std_logic;
   signal AC_ADR1 : std_logic;
   signal AC_GPIO0 : std_logic;
   signal AC_GPIO2 : std_logic;
   signal AC_GPIO3 : std_logic;
   signal AC_MCLK : std_logic;
   signal AC_SCK : std_logic;

   signal lr_stim  : std_logic_vector(63 downto 0) := x"FFFFFFFF00000000";
   signal d_stim   : std_logic_vector(63 downto 0) := x"4000000040000000";
   -- Clock period definitions
   constant clk_100_period : time := 10 ns;
BEGIN
   AC_SDA <= 'H';
   
	-- Instantiate the Unit Under Test (UUT)
   uut: adau1761_test PORT MAP (
          clk_100 => clk_100,
          AC_ADR0 => AC_ADR0,
          AC_ADR1 => AC_ADR1,
          AC_GPIO0 => AC_GPIO0,
          AC_GPIO1 => AC_GPIO1,
          AC_GPIO2 => AC_GPIO2,
          AC_GPIO3 => AC_GPIO3,
          AC_MCLK => AC_MCLK,
          AC_SCK => AC_SCK,
          AC_SDA => AC_SDA,
          sw=> "00000001"
        );

   -- Clock process definitions
   clk_100_process :process
   begin
		clk_100 <= '0';
		wait for clk_100_period/2;
		clk_100 <= '1';
		wait for clk_100_period/2;
   end process;
 
   AC_GPIO3 <= lr_stim(lr_stim'high);
   AC_GPIO1 <= d_stim(d_stim'high);


-- simulate the clocks generated by the codec chip.   
 i2s_clock : process
   begin
      AC_GPIO2 <= '1';
      wait for 1000000.0 ns /48/64/2;
      AC_GPIO2 <= '0';
      lr_stim <= lr_stim(lr_stim'high-1 downto 0) & lr_stim(lr_stim'high);
      d_stim  <= d_stim(d_stim'high-1 downto 0)   & d_stim(lr_stim'high);
      wait for 1000000.0 ns /48/64/2;
   end process;
   -- Stimulus process
   stim_proc: process
   begin		
      wait;
   end process;

END;
